grammar edu:umn:cs:melt:exts:ableC:allocation;

exports edu:umn:cs:melt:exts:ableC:allocation:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:allocation:abstractsyntax;