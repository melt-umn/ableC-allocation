grammar edu:umn:cs:melt:exts:ableC:allocation:concretesyntax;

imports edu:umn:cs:melt:ableC:concretesyntax;
imports edu:umn:cs:melt:ableC:abstractsyntax:host as ast;
imports edu:umn:cs:melt:ableC:abstractsyntax:construction as ast;
imports edu:umn:cs:melt:exts:ableC:allocation:abstractsyntax;

imports silver:langutil only ast;